module alu_top(
    input clk,
    input rst,
    input opcode,
    output funct
);

endmodule